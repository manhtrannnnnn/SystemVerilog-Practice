//----------------------------Last In First Out--------------------------------//
module lifo(
    input clk, 
    input [7:0] data_in, 
    input wr_en, rd_en,
    output empty, full,
    output logic [7:0] data_out
);



endmodule